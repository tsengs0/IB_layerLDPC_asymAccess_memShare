`ifndef __H_MEMSHARE_IBLUT_CONFIG
`define __H_MEMSHARE_IBLUT_CONFIG

//`define MEMSHARE_VN_IBRAM_BANK_INTERLEAVE

`endif // __H_MEMSHARE_IBLUT_CONFIG
