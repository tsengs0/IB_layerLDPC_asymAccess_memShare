parameter TRIAL0 = 3;
parameter TRIAL1 = 5;
parameter TRIAL2 = 9;
parameter TRIAL3 = 15;
parameter TRIAL4 = 17;
parameter TRIAL5 = 45;
parameter TRIAL6 = 51;
parameter TRIAL7 = 85;
parameter TRIAL8 = 153;
parameter TRIAL9 = 255;