module qsn_controller_len51 #(
	parameter [$clog2(51)-1:0] PERMUTATION_LENGTH = 51
) (
	output wire [5:0] left_sel,
	output wire [5:0] right_sel,
	output wire [49:0] merge_sel,
	input wire [5:0] shift_factor
//,	input wire rstn,
//	input wire sys_clk
);

	wire shifter_nonzero;
	assign shifter_nonzero = (|shift_factor[5:0]);

	assign left_sel[5:0] = (shifter_nonzero == 1'b1) ? shift_factor[5:0] : 0;
	assign right_sel[5:0] = (shifter_nonzero == 1'b1) ? 51-shift_factor[5:0] : 0;
	assign merge_sel[49:0] = f(shift_factor[5:0]);
	function [49:0] f(input [5:0] shift_in);
		case(shift_in[5:0])
			1	:	 f[49:0] = 50'b11111111111111111111111111111111111111111111111111;
			2	:	 f[49:0] = 50'b01111111111111111111111111111111111111111111111111;
			3	:	 f[49:0] = 50'b00111111111111111111111111111111111111111111111111;
			4	:	 f[49:0] = 50'b00011111111111111111111111111111111111111111111111;
			5	:	 f[49:0] = 50'b00001111111111111111111111111111111111111111111111;
			6	:	 f[49:0] = 50'b00000111111111111111111111111111111111111111111111;
			7	:	 f[49:0] = 50'b00000011111111111111111111111111111111111111111111;
			8	:	 f[49:0] = 50'b00000001111111111111111111111111111111111111111111;
			9	:	 f[49:0] = 50'b00000000111111111111111111111111111111111111111111;
			10	:	 f[49:0] = 50'b00000000011111111111111111111111111111111111111111;
			11	:	 f[49:0] = 50'b00000000001111111111111111111111111111111111111111;
			12	:	 f[49:0] = 50'b00000000000111111111111111111111111111111111111111;
			13	:	 f[49:0] = 50'b00000000000011111111111111111111111111111111111111;
			14	:	 f[49:0] = 50'b00000000000001111111111111111111111111111111111111;
			15	:	 f[49:0] = 50'b00000000000000111111111111111111111111111111111111;
			16	:	 f[49:0] = 50'b00000000000000011111111111111111111111111111111111;
			17	:	 f[49:0] = 50'b00000000000000001111111111111111111111111111111111;
			18	:	 f[49:0] = 50'b00000000000000000111111111111111111111111111111111;
			19	:	 f[49:0] = 50'b00000000000000000011111111111111111111111111111111;
			20	:	 f[49:0] = 50'b00000000000000000001111111111111111111111111111111;
			21	:	 f[49:0] = 50'b00000000000000000000111111111111111111111111111111;
			22	:	 f[49:0] = 50'b00000000000000000000011111111111111111111111111111;
			23	:	 f[49:0] = 50'b00000000000000000000001111111111111111111111111111;
			24	:	 f[49:0] = 50'b00000000000000000000000111111111111111111111111111;
			25	:	 f[49:0] = 50'b00000000000000000000000011111111111111111111111111;
			26	:	 f[49:0] = 50'b00000000000000000000000001111111111111111111111111;
			27	:	 f[49:0] = 50'b00000000000000000000000000111111111111111111111111;
			28	:	 f[49:0] = 50'b00000000000000000000000000011111111111111111111111;
			29	:	 f[49:0] = 50'b00000000000000000000000000001111111111111111111111;
			30	:	 f[49:0] = 50'b00000000000000000000000000000111111111111111111111;
			31	:	 f[49:0] = 50'b00000000000000000000000000000011111111111111111111;
			32	:	 f[49:0] = 50'b00000000000000000000000000000001111111111111111111;
			33	:	 f[49:0] = 50'b00000000000000000000000000000000111111111111111111;
			34	:	 f[49:0] = 50'b00000000000000000000000000000000011111111111111111;
			35	:	 f[49:0] = 50'b00000000000000000000000000000000001111111111111111;
			36	:	 f[49:0] = 50'b00000000000000000000000000000000000111111111111111;
			37	:	 f[49:0] = 50'b00000000000000000000000000000000000011111111111111;
			38	:	 f[49:0] = 50'b00000000000000000000000000000000000001111111111111;
			39	:	 f[49:0] = 50'b00000000000000000000000000000000000000111111111111;
			40	:	 f[49:0] = 50'b00000000000000000000000000000000000000011111111111;
			41	:	 f[49:0] = 50'b00000000000000000000000000000000000000001111111111;
			42	:	 f[49:0] = 50'b00000000000000000000000000000000000000000111111111;
			43	:	 f[49:0] = 50'b00000000000000000000000000000000000000000011111111;
			44	:	 f[49:0] = 50'b00000000000000000000000000000000000000000001111111;
			45	:	 f[49:0] = 50'b00000000000000000000000000000000000000000000111111;
			46	:	 f[49:0] = 50'b00000000000000000000000000000000000000000000011111;
			47	:	 f[49:0] = 50'b00000000000000000000000000000000000000000000001111;
			48	:	 f[49:0] = 50'b00000000000000000000000000000000000000000000000111;
			49	:	 f[49:0] = 50'b00000000000000000000000000000000000000000000000011;
			50	:	 f[49:0] = 50'b00000000000000000000000000000000000000000000000001;
			default	:	f[49:0] = 0;
		endcase // shift_factor
	endfunction
endmodule