class scu_memShare_tb_class;

task dirver;

endtask

endclass
