package scu_memShare_tb_config_pkg;

localparam TB_CLK_DELAY = 0; // Delay from the starting point
localparam TB_CLK_PERIOD = 10;
localparam logic TB_CLK_INITAL_LEVEL = 1'b0;
endpackage: scu_memShare_tb_config_pkg
