`ifndef __GLOBAL_DEBUG_H
`define __GLOBAL_DEBUG_H

//`define TB_DEBUG

`endif // __GLOBAL_DEBUG_H
